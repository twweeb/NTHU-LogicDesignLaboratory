`timescale 1ns / 1ps

module Ground (
    input wire clk,
    input wire [8:0] row_addr,
    input wire [9:0] col_addr,
    output reg [9:0] ground_position,
    input wire game_status,
    input wire fresh,
    output reg [3:0] speed,
    output reg px
    );
    reg [159:0] pattern [7:0];

    always @(negedge fresh) begin
        if (game_status) begin
            ground_position<=(ground_position+speed)%10'd160;//move the ground
        end
    end

    always @(posedge clk) //begin
    begin
        if (row_addr>=10'd400 && row_addr<10'd408) begin
            px <= pattern[row_addr-10'd400][(col_addr+ground_position)%10'd160];
        end else begin
            px <= 1'b0;
        end
        if (game_status==1'b0) begin
            speed<=4'd6;
            pattern[0]<=160'b1010111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111;
            pattern[1]<=160'b0101000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000;
            pattern[2]<=160'b0000000000011100000000000000000000000011100000000000000000000000000000000000000000000001100000000000000000000001110000000000000000000000000000000000000000000000;
            pattern[3]<=160'b0000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000;
            pattern[4]<=160'b0000000000010000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000;
            pattern[5]<=160'b0000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000;
            pattern[6]<=160'b0000000010000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000111000000000000000000000000000;
            pattern[7]<=160'b0000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
        end
    end
    
    initial begin
        ground_position<=10'b0;
    end
    

endmodule

