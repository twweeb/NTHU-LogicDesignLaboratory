`timescale 1ns / 1ps

module Jump (
    input wire fresh,
    input wire clk,
    input wire jump,
    input wire RESET,
    input wire START,
    input wire [8:0] row_addr,
    input wire [9:0] col_addr,
    output reg px, // Display
    input wire game_status
    );
    
    reg [11:0] jump_time;
    wire [11:0] height;
    reg [0:82] run [0:49];
    reg is_jumping;

    reg [3:0] counter;

    //height is only associated with the value of jump_time
    assign height = (jump_time*12'd40 - jump_time*jump_time) / 2'd2;

    // every frame
    always @(negedge fresh) begin
        counter<=counter+1;
        if (game_status) begin
            if (jump && is_jumping==1'b0) begin
               is_jumping<=1'b1;//begin to jump
            end
            if (is_jumping) begin
                if (jump_time>=12'd40) begin//reset jump operation
                    jump_time<=12'b0;
                    is_jumping<=1'b0;
                end else begin
                    jump_time<=jump_time+1'b1;//add jump_time
                end
            end
        end else begin //if pausing
            if (RESET || START) begin
                jump_time<=12'b0;
                is_jumping<=1'b0;
                counter<=4'b0;
            end
        end
        
    end

    always @(posedge clk) begin
        //body part is based on row_addr and col_addr
        if (row_addr >= 10'd402 - height - 10'd50 && row_addr < 10'd402 - height && col_addr>=10'd80 && col_addr<10'd162) begin
            px <= run[row_addr+height-10'd352][col_addr-12'd80];
        end else begin
            px <= 1'b0;
        end
    end

    always @(posedge RESET) begin
        //use ram to store the pattern of dinosaur (row 88, col 82)
        run[0] <=82'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        run[1] <=82'b0000000000000000000000000000000000000000000000000000000000000000011111000001000000;
        run[2] <=82'b0000000000000000000000000000000000000000000000000000000000000111111111111111111000;
        run[3] <=82'b0000000000000000000000000000000000000000000000000000000000011111111101111111111100;
        run[4] <=82'b0000000000000000000000000000000000000000000000000000000000111111111101111111111110;
        run[5] <=82'b0000000000000000000000000000000000000000000000000000000001111111111111111111111110;
        run[6] <=82'b0000000000000000000000000000000000000000000000000000000011111111111111111111111110;
        run[7] <=82'b0000000000000000000000000000000000000000000000000000000111111111011111111010010000;
        run[8] <=82'b0000000000000000000000000000000000000000111111111000011111111111111111000000010000;
        run[9] <=82'b0000000000000000000000000000011111111111111111111111111111111111111110000000000000;
        run[10]<=82'b0000000000000000000000000011111111111111111111111111111111111111111110000000000000;
        run[11]<=82'b0000000000000000000000001111111111111111111111111111111111111111111111000000000000;
        run[12]<=82'b0000000000000000000000011111111111111111111111111111111111111111111111100000000000;
        run[13]<=82'b0000000000000000000001111111111111111111111111111111111111111111111111110000000000;
        run[14]<=82'b0000000000000000001111111111111111111111111111111111111111111111111111111100000000;
        run[15]<=82'b0000000000000001111111111111111111111111111111111111111111111111111111111110000000;
        run[16]<=82'b0000000000111111111111111111111111111111111111111111111111111111000011111111110000;
        run[17]<=82'b0000000111111111111111111111111111111111111111111111111111111100000000001111110000;
        run[18]<=82'b0000011111111111111111111111111111111111111111111111111111111000000000000011110000;
        run[19]<=82'b0000111111111111111111111111100111111111111111111111111111000000000000000000000000;
        run[20]<=82'b0001111111111111111111111111110011111111111111111111111110000000000000000000000000;
        run[21]<=82'b0011111111111111111111111111111101111111111111111111111100000000000000000000000000;
        run[22]<=82'b0111111111111111111111111111111110111111111111111111111000000000000000000000000000;
        run[23]<=82'b0111111111111111111111111111111111111111111111111111111000000000000000000000000000;
        run[24]<=82'b0111100000000000000111111011111111111111111111111111111000000000000000000000000000;
        run[25]<=82'b1111000000000000000000111110111111111111111111111111011110001000000000000000000000;
        run[26]<=82'b0111000000000000000000011111011111111111111110000010001111110000000000000000000000;
        run[27]<=82'b0111000000000000000000000000111111111111110000000001000000001000000000000000000000;
        run[28]<=82'b0111000000000000000000000000001111111100000000000000000000000000000000000000000000;
        run[29]<=82'b0011110000000000000000000000001110111100000000000000000000000000000000000000000000;
        run[30]<=82'b0001111000000000000000000000111111111000000000000000000000000000000000000000000000;
        run[31]<=82'b0000011110000000000000000001111111111000000000000000000000000000000000000000000000;
        run[32]<=82'b0000000011000000000000000011111111111000000000000000000000000000000000000000000000;
        run[33]<=82'b0000000000110000000000111111111111110000000000000000000000000000000000000000000000;
        run[34]<=82'b0000000000010000000001111111111111000000000000000000000000000000000000000000000000;
        run[35]<=82'b0000000000010000000011111111111110000000000000000000000000000000000000000000000000;
        run[36]<=82'b0000000000010000000111111000111100000000000000000000000000000000000000000000000000;
        run[37]<=82'b0000000000000000000111110001111100000000000000000000000000000000000000000000000000;
        run[38]<=82'b0000000000000000000111100001111000000000000000000000000000000000000000000000000000;
        run[39]<=82'b0000000000000000001111100000111000000000000000000000000000000000000000000000000000;
        run[40]<=82'b0000000000000000001111100000111000000000000000000000000000000000000000000000000000;
        run[41]<=82'b0000000000000000001111100000111100000000000000000000000000000000000000000000000000;
        run[42]<=82'b0000000000000000001111100000011100000000000000000000000000000000000000000000000000;
        run[43]<=82'b0000000000000000000111100000011110000000000000000000000000000000000000000000000000;
        run[44]<=82'b0000000000000000000111110000011111000000000000000000000000000000000000000000000000;
        run[45]<=82'b0000000000000000000011111100011111100000000000000000000000000000000000000000000000;
        run[46]<=82'b0000000000000000000000000000011111111111000000000000000000000000000000000000000000;
        run[47]<=82'b0000000000000000000000000000011111111110000000000000000000000000000000000000000000;
        run[48]<=82'b0000000000000000000000000000001100011000000000000000000000000000000000000000000000;
        run[49]<=82'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      end
    
 
    
endmodule
