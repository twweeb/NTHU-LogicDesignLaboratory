`define s1  32'd524 // C sharp
`define s2  32'd588 // D sharp
`define s3  32'd660 // E sharp
`define s4  32'd698 // F sharp
`define s5  32'd784 // G sharp
`define s6  32'd880 // A sharp
`define s7  32'd988 // B sharp
`define n1   32'd262 // C
`define n2   32'd294 // E
`define n3   32'd330 // D
`define n4   32'd349 // F
`define n5   32'd392 // G
`define n6   32'd440 // A
`define n7   32'd494 // B
`define sil   32'd50000000 // slience

//Frere Jacques
module music (
    input [11:0] ibeatNum,
    input en,
    output reg [31:0] toneL,
    output reg [31:0] toneR
);

    always @* begin
        if(en == 0) begin
            case(ibeatNum)
                12'd0: toneR = `s1;    12'd1: toneR = `s1;    12'd2: toneR = `s1;    12'd3: toneR = `s1;    12'd4: toneR = `s1;    12'd5: toneR = `s1;    12'd6: toneR = `s1;    12'd7: toneR = `s1;    12'd8: toneR = `s1;    12'd9: toneR = `s1;    12'd10: toneR = `s1;    12'd11: toneR = `s1;    12'd12: toneR = `s1;    12'd13: toneR = `s1;    12'd14: toneR = `s1;    12'd15: toneR = `sil;    12'd16: toneR = `s2;    12'd17: toneR = `s2;    12'd18: toneR = `s2;    12'd19: toneR = `s2;    12'd20: toneR = `s2;    12'd21: toneR = `s2;    12'd22: toneR = `s2;    12'd23: toneR = `s2;    12'd24: toneR = `s2;    12'd25: toneR = `s2;    12'd26: toneR = `s2;    12'd27: toneR = `s2;    12'd28: toneR = `s2;    12'd29: toneR = `s2;    12'd30: toneR = `s2;    12'd31: toneR = `sil;    12'd32: toneR = `s3;    12'd33: toneR = `s3;    12'd34: toneR = `s3;    12'd35: toneR = `s3;    12'd36: toneR = `s3;    12'd37: toneR = `s3;    12'd38: toneR = `s3;    12'd39: toneR = `s3;    12'd40: toneR = `s3;    12'd41: toneR = `s3;    12'd42: toneR = `s3;    12'd43: toneR = `s3;    12'd44: toneR = `s3;    12'd45: toneR = `s3;    12'd46: toneR = `s3;    12'd47: toneR = `sil;    12'd48: toneR = `s1;    12'd49: toneR = `s1;    12'd50: toneR = `s1;    12'd51: toneR = `s1;    12'd52: toneR = `s1;    12'd53: toneR = `s1;    12'd54: toneR = `s1;    12'd55: toneR = `s1;    12'd56: toneR = `s1;    12'd57: toneR = `s1;    12'd58: toneR = `s1;    12'd59: toneR = `s1;    12'd60: toneR = `s1;    12'd61: toneR = `s1;    12'd62: toneR = `s1;    12'd63: toneR = `sil;
                12'd64: toneR = `s1;    12'd65: toneR = `s1;    12'd66: toneR = `s1;    12'd67: toneR = `s1;    12'd68: toneR = `s1;    12'd69: toneR = `s1;    12'd70: toneR = `s1;    12'd71: toneR = `s1;    12'd72: toneR = `s1;    12'd73: toneR = `s1;    12'd74: toneR = `s1;    12'd75: toneR = `s1;    12'd76: toneR = `s1;    12'd77: toneR = `s1;    12'd78: toneR = `s1;    12'd79: toneR = `sil;    12'd80: toneR = `s2;    12'd81: toneR = `s2;    12'd82: toneR = `s2;    12'd83: toneR = `s2;    12'd84: toneR = `s2;    12'd85: toneR = `s2;    12'd86: toneR = `s2;    12'd87: toneR = `s2;    12'd88: toneR = `s2;    12'd89: toneR = `s2;    12'd90: toneR = `s2;    12'd91: toneR = `s2;    12'd92: toneR = `s2;    12'd93: toneR = `s2;    12'd94: toneR = `s2;    12'd95: toneR = `sil;    12'd96: toneR = `s3;    12'd97: toneR = `s3;    12'd98: toneR = `s3;    12'd99: toneR = `s3;    12'd100: toneR = `s3;    12'd101: toneR = `s3;    12'd102: toneR = `s3;    12'd103: toneR = `s3;    12'd104: toneR = `s3;    12'd105: toneR = `s3;    12'd106: toneR = `s3;    12'd107: toneR = `s3;    12'd108: toneR = `s3;    12'd109: toneR = `s3;    12'd110: toneR = `s3;    12'd111: toneR = `sil;    12'd112: toneR = `s1;    12'd113: toneR = `s1;    12'd114: toneR = `s1;    12'd115: toneR = `s1;    12'd116: toneR = `s1;    12'd117: toneR = `s1;    12'd118: toneR = `s1;    12'd119: toneR = `s1;    12'd120: toneR = `s1;    12'd121: toneR = `s1;    12'd122: toneR = `s1;    12'd123: toneR = `s1;    12'd124: toneR = `s1;    12'd125: toneR = `s1;    12'd126: toneR = `s1;    12'd127: toneR = `sil;
                12'd128: toneR = `s3;    12'd129: toneR = `s3;    12'd130: toneR = `s3;    12'd131: toneR = `s3;    12'd132: toneR = `s3;    12'd133: toneR = `s3;    12'd134: toneR = `s3;    12'd135: toneR = `s3;    12'd136: toneR = `s3;    12'd137: toneR = `s3;    12'd138: toneR = `s3;    12'd139: toneR = `s3;    12'd140: toneR = `s3;    12'd141: toneR = `s3;    12'd142: toneR = `s3;    12'd143: toneR = `sil;    12'd144: toneR = `s4;    12'd145: toneR = `s4;    12'd146: toneR = `s4;    12'd147: toneR = `s4;    12'd148: toneR = `s4;    12'd149: toneR = `s4;    12'd150: toneR = `s4;    12'd151: toneR = `s4;    12'd152: toneR = `s4;    12'd153: toneR = `s4;    12'd154: toneR = `s4;    12'd155: toneR = `s4;    12'd156: toneR = `s4;    12'd157: toneR = `s4;    12'd158: toneR = `s4;    12'd159: toneR = `sil;    12'd160: toneR = `s5;    12'd161: toneR = `s5;    12'd162: toneR = `s5;    12'd163: toneR = `s5;    12'd164: toneR = `s5;    12'd165: toneR = `s5;    12'd166: toneR = `s5;    12'd167: toneR = `s5;    12'd168: toneR = `s5;    12'd169: toneR = `s5;    12'd170: toneR = `s5;    12'd171: toneR = `s5;    12'd172: toneR = `s5;    12'd173: toneR = `s5;    12'd174: toneR = `s5;    12'd175: toneR = `s5;    12'd176: toneR = `s5;    12'd177: toneR = `s5;    12'd178: toneR = `s5;    12'd179: toneR = `s5;    12'd180: toneR = `s5;    12'd181: toneR = `s5;    12'd182: toneR = `s5;    12'd183: toneR = `s5;    12'd184: toneR = `s5;    12'd185: toneR = `s5;    12'd186: toneR = `s5;    12'd187: toneR = `s5;    12'd188: toneR = `s5;    12'd189: toneR = `s5;    12'd190: toneR = `s5;    12'd191: toneR = `sil;
                12'd192: toneR = `s3;    12'd193: toneR = `s3;    12'd194: toneR = `s3;    12'd195: toneR = `s3;    12'd196: toneR = `s3;    12'd197: toneR = `s3;    12'd198: toneR = `s3;    12'd199: toneR = `s3;    12'd200: toneR = `s3;    12'd201: toneR = `s3;    12'd202: toneR = `s3;    12'd203: toneR = `s3;    12'd204: toneR = `s3;    12'd205: toneR = `s3;    12'd206: toneR = `s3;    12'd207: toneR = `sil;    12'd208: toneR = `s4;    12'd209: toneR = `s4;    12'd210: toneR = `s4;    12'd211: toneR = `s4;    12'd212: toneR = `s4;    12'd213: toneR = `s4;    12'd214: toneR = `s4;    12'd215: toneR = `s4;    12'd216: toneR = `s4;    12'd217: toneR = `s4;    12'd218: toneR = `s4;    12'd219: toneR = `s4;    12'd220: toneR = `s4;    12'd221: toneR = `s4;    12'd222: toneR = `s4;    12'd223: toneR = `sil;    12'd224: toneR = `s5;    12'd225: toneR = `s5;    12'd226: toneR = `s5;    12'd227: toneR = `s5;    12'd228: toneR = `s5;    12'd229: toneR = `s5;    12'd230: toneR = `s5;    12'd231: toneR = `s5;    12'd232: toneR = `s5;    12'd233: toneR = `s5;    12'd234: toneR = `s5;    12'd235: toneR = `s5;    12'd236: toneR = `s5;    12'd237: toneR = `s5;    12'd238: toneR = `s5;    12'd239: toneR = `s5;    12'd240: toneR = `s5;    12'd241: toneR = `s5;    12'd242: toneR = `s5;    12'd243: toneR = `s5;    12'd244: toneR = `s5;    12'd245: toneR = `s5;    12'd246: toneR = `s5;    12'd247: toneR = `s5;    12'd248: toneR = `s5;    12'd249: toneR = `s5;    12'd250: toneR = `s5;    12'd251: toneR = `s5;    12'd252: toneR = `s5;    12'd253: toneR = `s5;    12'd254: toneR = `s5;    12'd255: toneR = `sil;
                12'd256: toneR = `s5;    12'd257: toneR = `s5;    12'd258: toneR = `s5;    12'd259: toneR = `s5;    12'd260: toneR = `s5;    12'd261: toneR = `s5;    12'd262: toneR = `s5;    12'd263: toneR = `s5;    12'd264: toneR = `s6;    12'd265: toneR = `s6;    12'd266: toneR = `s6;    12'd267: toneR = `s6;    12'd268: toneR = `s6;    12'd269: toneR = `s6;    12'd270: toneR = `s6;    12'd271: toneR = `s6;    12'd272: toneR = `s5;    12'd273: toneR = `s5;    12'd274: toneR = `s5;    12'd275: toneR = `s5;    12'd276: toneR = `s5;    12'd277: toneR = `s5;    12'd278: toneR = `s5;    12'd279: toneR = `s5;    12'd280: toneR = `s4;    12'd281: toneR = `s4;    12'd282: toneR = `s4;    12'd283: toneR = `s4;    12'd284: toneR = `s4;    12'd285: toneR = `s4;    12'd286: toneR = `s4;    12'd287: toneR = `sil;    12'd288: toneR = `s3;    12'd289: toneR = `s3;    12'd290: toneR = `s3;    12'd291: toneR = `s3;    12'd292: toneR = `s3;    12'd293: toneR = `s3;    12'd294: toneR = `s3;    12'd295: toneR = `s3;    12'd296: toneR = `s3;    12'd297: toneR = `s3;    12'd298: toneR = `s3;    12'd299: toneR = `s3;    12'd300: toneR = `s3;    12'd301: toneR = `s3;    12'd302: toneR = `s3;    12'd303: toneR = `sil;    12'd304: toneR = `s1;    12'd305: toneR = `s1;    12'd306: toneR = `s1;    12'd307: toneR = `s1;    12'd308: toneR = `s1;    12'd309: toneR = `s1;    12'd310: toneR = `s1;    12'd311: toneR = `s1;    12'd312: toneR = `s1;    12'd313: toneR = `s1;    12'd314: toneR = `s1;    12'd315: toneR = `s1;    12'd316: toneR = `s1;    12'd317: toneR = `s1;    12'd318: toneR = `s1;    12'd319: toneR = `sil;
                12'd320: toneR = `s5;    12'd321: toneR = `s5;    12'd322: toneR = `s5;    12'd323: toneR = `s5;    12'd324: toneR = `s5;    12'd325: toneR = `s5;    12'd326: toneR = `s5;    12'd327: toneR = `s5;    12'd328: toneR = `s6;    12'd329: toneR = `s6;    12'd330: toneR = `s6;    12'd331: toneR = `s6;    12'd332: toneR = `s6;    12'd333: toneR = `s6;    12'd334: toneR = `s6;    12'd335: toneR = `s6;    12'd336: toneR = `s5;    12'd337: toneR = `s5;    12'd338: toneR = `s5;    12'd339: toneR = `s5;    12'd340: toneR = `s5;    12'd341: toneR = `s5;    12'd342: toneR = `s5;    12'd343: toneR = `s5;    12'd344: toneR = `s4;    12'd345: toneR = `s4;    12'd346: toneR = `s4;    12'd347: toneR = `s4;    12'd348: toneR = `s4;    12'd349: toneR = `s4;    12'd350: toneR = `s4;    12'd351: toneR = `sil;    12'd352: toneR = `s3;    12'd353: toneR = `s3;    12'd354: toneR = `s3;    12'd355: toneR = `s3;    12'd356: toneR = `s3;    12'd357: toneR = `s3;    12'd358: toneR = `s3;    12'd359: toneR = `s3;    12'd360: toneR = `s3;    12'd361: toneR = `s3;    12'd362: toneR = `s3;    12'd363: toneR = `s3;    12'd364: toneR = `s3;    12'd365: toneR = `s3;    12'd366: toneR = `s3;    12'd367: toneR = `sil;    12'd368: toneR = `s1;    12'd369: toneR = `s1;    12'd370: toneR = `s1;    12'd371: toneR = `s1;    12'd372: toneR = `s1;    12'd373: toneR = `s1;    12'd374: toneR = `s1;    12'd375: toneR = `s1;    12'd376: toneR = `s1;    12'd377: toneR = `s1;    12'd378: toneR = `s1;    12'd379: toneR = `s1;    12'd380: toneR = `s1;    12'd381: toneR = `s1;    12'd382: toneR = `s1;    12'd383: toneR = `sil;
                12'd384: toneR = `s1;    12'd385: toneR = `s1;    12'd386: toneR = `s1;    12'd387: toneR = `s1;    12'd388: toneR = `s1;    12'd389: toneR = `s1;    12'd390: toneR = `s1;    12'd391: toneR = `s1;    12'd392: toneR = `s1;    12'd393: toneR = `s1;    12'd394: toneR = `s1;    12'd395: toneR = `s1;    12'd396: toneR = `s1;    12'd397: toneR = `s1;    12'd398: toneR = `s1;    12'd399: toneR = `sil;    12'd400: toneR = `n5;    12'd401: toneR = `n5;    12'd402: toneR = `n5;    12'd403: toneR = `n5;    12'd404: toneR = `n5;    12'd405: toneR = `n5;    12'd406: toneR = `n5;    12'd407: toneR = `n5;    12'd408: toneR = `n5;    12'd409: toneR = `n5;    12'd410: toneR = `n5;    12'd411: toneR = `n5;    12'd412: toneR = `n5;    12'd413: toneR = `n5;    12'd414: toneR = `n5;    12'd415: toneR = `sil;    12'd416: toneR = `s1;    12'd417: toneR = `s1;    12'd418: toneR = `s1;    12'd419: toneR = `s1;    12'd420: toneR = `s1;    12'd421: toneR = `s1;    12'd422: toneR = `s1;    12'd423: toneR = `s1;    12'd424: toneR = `s1;    12'd425: toneR = `s1;    12'd426: toneR = `s1;    12'd427: toneR = `s1;    12'd428: toneR = `s1;    12'd429: toneR = `s1;    12'd430: toneR = `s1;    12'd431: toneR = `s1;    12'd432: toneR = `s1;    12'd433: toneR = `s1;    12'd434: toneR = `s1;    12'd435: toneR = `s1;    12'd436: toneR = `s1;    12'd437: toneR = `s1;    12'd438: toneR = `s1;    12'd439: toneR = `s1;    12'd440: toneR = `s1;    12'd441: toneR = `s1;    12'd442: toneR = `s1;    12'd443: toneR = `s1;    12'd444: toneR = `s1;    12'd445: toneR = `s1;    12'd446: toneR = `s1;    12'd447: toneR = `sil;
                12'd448: toneR = `s1;    12'd449: toneR = `s1;    12'd450: toneR = `s1;    12'd451: toneR = `s1;    12'd452: toneR = `s1;    12'd453: toneR = `s1;    12'd454: toneR = `s1;    12'd455: toneR = `s1;    12'd456: toneR = `s1;    12'd457: toneR = `s1;    12'd458: toneR = `s1;    12'd459: toneR = `s1;    12'd460: toneR = `s1;    12'd461: toneR = `s1;    12'd462: toneR = `s1;    12'd463: toneR = `sil;    12'd464: toneR = `n5;    12'd465: toneR = `n5;    12'd466: toneR = `n5;    12'd467: toneR = `n5;    12'd468: toneR = `n5;    12'd469: toneR = `n5;    12'd470: toneR = `n5;    12'd471: toneR = `n5;    12'd472: toneR = `n5;    12'd473: toneR = `n5;    12'd474: toneR = `n5;    12'd475: toneR = `n5;    12'd476: toneR = `n5;    12'd477: toneR = `n5;    12'd478: toneR = `n5;    12'd479: toneR = `sil;    12'd480: toneR = `s1;    12'd481: toneR = `s1;    12'd482: toneR = `s1;    12'd483: toneR = `s1;    12'd484: toneR = `s1;    12'd485: toneR = `s1;    12'd486: toneR = `s1;    12'd487: toneR = `s1;    12'd488: toneR = `s1;    12'd489: toneR = `s1;    12'd490: toneR = `s1;    12'd491: toneR = `s1;    12'd492: toneR = `s1;    12'd493: toneR = `s1;    12'd494: toneR = `s1;    12'd495: toneR = `s1;    12'd496: toneR = `s1;    12'd497: toneR = `s1;    12'd498: toneR = `s1;    12'd499: toneR = `s1;    12'd500: toneR = `s1;    12'd501: toneR = `s1;    12'd502: toneR = `s1;    12'd503: toneR = `s1;    12'd504: toneR = `s1;    12'd505: toneR = `s1;    12'd506: toneR = `s1;    12'd507: toneR = `s1;    12'd508: toneR = `s1;    12'd509: toneR = `s1;    12'd510: toneR = `s1;    12'd511: toneR = `sil;
                default : toneR = `sil;
            endcase
        end else begin
            toneR = `sil;
        end
    end

    always @(*) begin
        if(en==0)begin
            case(ibeatNum)
                12'd0: toneL = `s1;    12'd1: toneL = `s1;    12'd2: toneL = `s1;    12'd3: toneL = `s1;    12'd4: toneL = `s1;    12'd5: toneL = `s1;    12'd6: toneL = `s1;    12'd7: toneL = `s1;    12'd8: toneL = `s1;    12'd9: toneL = `s1;    12'd10: toneL = `s1;    12'd11: toneL = `s1;    12'd12: toneL = `s1;    12'd13: toneL = `s1;    12'd14: toneL = `s1;    12'd15: toneL = `s1;    12'd16: toneL = `s1;    12'd17: toneL = `s1;    12'd18: toneL = `s1;    12'd19: toneL = `s1;    12'd20: toneL = `s1;    12'd21: toneL = `s1;    12'd22: toneL = `s1;    12'd23: toneL = `s1;    12'd24: toneL = `s1;    12'd25: toneL = `s1;    12'd26: toneL = `s1;    12'd27: toneL = `s1;    12'd28: toneL = `s1;    12'd29: toneL = `s1;    12'd30: toneL = `s1;    12'd31: toneL = `sil;    12'd32: toneL = `n5;    12'd33: toneL = `n5;    12'd34: toneL = `n5;    12'd35: toneL = `n5;    12'd36: toneL = `n5;    12'd37: toneL = `n5;    12'd38: toneL = `n5;    12'd39: toneL = `n5;    12'd40: toneL = `n5;    12'd41: toneL = `n5;    12'd42: toneL = `n5;    12'd43: toneL = `n5;    12'd44: toneL = `n5;    12'd45: toneL = `n5;    12'd46: toneL = `n5;    12'd47: toneL = `n5;    12'd48: toneL = `n5;    12'd49: toneL = `n5;    12'd50: toneL = `n5;    12'd51: toneL = `n5;    12'd52: toneL = `n5;    12'd53: toneL = `n5;    12'd54: toneL = `n5;    12'd55: toneL = `n5;    12'd56: toneL = `n5;    12'd57: toneL = `n5;    12'd58: toneL = `n5;    12'd59: toneL = `n5;    12'd60: toneL = `n5;    12'd61: toneL = `n5;    12'd62: toneL = `n5;    12'd63: toneL = `sil;
                12'd64: toneL = `s1;    12'd65: toneL = `s1;    12'd66: toneL = `s1;    12'd67: toneL = `s1;    12'd68: toneL = `s1;    12'd69: toneL = `s1;    12'd70: toneL = `s1;    12'd71: toneL = `s1;    12'd72: toneL = `s1;    12'd73: toneL = `s1;    12'd74: toneL = `s1;    12'd75: toneL = `s1;    12'd76: toneL = `s1;    12'd77: toneL = `s1;    12'd78: toneL = `s1;    12'd79: toneL = `s1;    12'd80: toneL = `s1;    12'd81: toneL = `s1;    12'd82: toneL = `s1;    12'd83: toneL = `s1;    12'd84: toneL = `s1;    12'd85: toneL = `s1;    12'd86: toneL = `s1;    12'd87: toneL = `s1;    12'd88: toneL = `s1;    12'd89: toneL = `s1;    12'd90: toneL = `s1;    12'd91: toneL = `s1;    12'd92: toneL = `s1;    12'd93: toneL = `s1;    12'd94: toneL = `s1;    12'd95: toneL = `sil;    12'd96: toneL = `n5;    12'd97: toneL = `n5;    12'd98: toneL = `n5;    12'd99: toneL = `n5;    12'd100: toneL = `n5;    12'd101: toneL = `n5;    12'd102: toneL = `n5;    12'd103: toneL = `n5;    12'd104: toneL = `n5;    12'd105: toneL = `n5;    12'd106: toneL = `n5;    12'd107: toneL = `n5;    12'd108: toneL = `n5;    12'd109: toneL = `n5;    12'd110: toneL = `n5;    12'd111: toneL = `n5;    12'd112: toneL = `n5;    12'd113: toneL = `n5;    12'd114: toneL = `n5;    12'd115: toneL = `n5;    12'd116: toneL = `n5;    12'd117: toneL = `n5;    12'd118: toneL = `n5;    12'd119: toneL = `n5;    12'd120: toneL = `n5;    12'd121: toneL = `n5;    12'd122: toneL = `n5;    12'd123: toneL = `n5;    12'd124: toneL = `n5;    12'd125: toneL = `n5;    12'd126: toneL = `n5;    12'd127: toneL = `sil;
                12'd128: toneL = `n1;    12'd129: toneL = `n1;    12'd130: toneL = `n1;    12'd131: toneL = `n1;    12'd132: toneL = `n1;    12'd133: toneL = `n1;    12'd134: toneL = `n1;    12'd135: toneL = `n1;    12'd136: toneL = `n1;    12'd137: toneL = `n1;    12'd138: toneL = `n1;    12'd139: toneL = `n1;    12'd140: toneL = `n1;    12'd141: toneL = `n1;    12'd142: toneL = `n1;    12'd143: toneL = `sil;    12'd144: toneL = `n2;    12'd145: toneL = `n2;    12'd146: toneL = `n2;    12'd147: toneL = `n2;    12'd148: toneL = `n2;    12'd149: toneL = `n2;    12'd150: toneL = `n2;    12'd151: toneL = `n2;    12'd152: toneL = `n2;    12'd153: toneL = `n2;    12'd154: toneL = `n2;    12'd155: toneL = `n2;    12'd156: toneL = `n2;    12'd157: toneL = `n2;    12'd158: toneL = `n2;    12'd159: toneL = `sil;    12'd160: toneL = `n3;    12'd161: toneL = `n3;    12'd162: toneL = `n3;    12'd163: toneL = `n3;    12'd164: toneL = `n3;    12'd165: toneL = `n3;    12'd166: toneL = `n3;    12'd167: toneL = `n3;    12'd168: toneL = `n3;    12'd169: toneL = `n3;    12'd170: toneL = `n3;    12'd171: toneL = `n3;    12'd172: toneL = `n3;    12'd173: toneL = `n3;    12'd174: toneL = `n3;    12'd175: toneL = `n3;    12'd176: toneL = `n3;    12'd177: toneL = `n3;    12'd178: toneL = `n3;    12'd179: toneL = `n3;    12'd180: toneL = `n3;    12'd181: toneL = `n3;    12'd182: toneL = `n3;    12'd183: toneL = `n3;    12'd184: toneL = `n3;    12'd185: toneL = `n3;    12'd186: toneL = `n3;    12'd187: toneL = `n3;    12'd188: toneL = `n3;    12'd189: toneL = `n3;    12'd190: toneL = `n3;    12'd191: toneL = `sil;
                12'd192: toneL = `n1;    12'd193: toneL = `n1;    12'd194: toneL = `n1;    12'd195: toneL = `n1;    12'd196: toneL = `n1;    12'd197: toneL = `n1;    12'd198: toneL = `n1;    12'd199: toneL = `n1;    12'd200: toneL = `n1;    12'd201: toneL = `n1;    12'd202: toneL = `n1;    12'd203: toneL = `n1;    12'd204: toneL = `n1;    12'd205: toneL = `n1;    12'd206: toneL = `n1;    12'd207: toneL = `sil;    12'd208: toneL = `n2;    12'd209: toneL = `n2;    12'd210: toneL = `n2;    12'd211: toneL = `n2;    12'd212: toneL = `n2;    12'd213: toneL = `n2;    12'd214: toneL = `n2;    12'd215: toneL = `n2;    12'd216: toneL = `n2;    12'd217: toneL = `n2;    12'd218: toneL = `n2;    12'd219: toneL = `n2;    12'd220: toneL = `n2;    12'd221: toneL = `n2;    12'd222: toneL = `n2;    12'd223: toneL = `sil;    12'd224: toneL = `n3;    12'd225: toneL = `n3;    12'd226: toneL = `n3;    12'd227: toneL = `n3;    12'd228: toneL = `n3;    12'd229: toneL = `n3;    12'd230: toneL = `n3;    12'd231: toneL = `n3;    12'd232: toneL = `n3;    12'd233: toneL = `n3;    12'd234: toneL = `n3;    12'd235: toneL = `n3;    12'd236: toneL = `n3;    12'd237: toneL = `n3;    12'd238: toneL = `n3;    12'd239: toneL = `n3;    12'd240: toneL = `n3;    12'd241: toneL = `n3;    12'd242: toneL = `n3;    12'd243: toneL = `n3;    12'd244: toneL = `n3;    12'd245: toneL = `n3;    12'd246: toneL = `n3;    12'd247: toneL = `n3;    12'd248: toneL = `n3;    12'd249: toneL = `n3;    12'd250: toneL = `n3;    12'd251: toneL = `n3;    12'd252: toneL = `n3;    12'd253: toneL = `n3;    12'd254: toneL = `n3;    12'd255: toneL = `sil;
                12'd256: toneL = `n3;    12'd257: toneL = `n3;    12'd258: toneL = `n3;    12'd259: toneL = `n3;    12'd260: toneL = `n3;    12'd261: toneL = `n3;    12'd262: toneL = `n3;    12'd263: toneL = `n3;    12'd264: toneL = `n3;    12'd265: toneL = `n3;    12'd266: toneL = `n3;    12'd267: toneL = `n3;    12'd268: toneL = `n3;    12'd269: toneL = `n3;    12'd270: toneL = `n3;    12'd271: toneL = `sil;    12'd272: toneL = `n4;    12'd273: toneL = `n4;    12'd274: toneL = `n4;    12'd275: toneL = `n4;    12'd276: toneL = `n4;    12'd277: toneL = `n4;    12'd278: toneL = `n4;    12'd279: toneL = `n4;    12'd280: toneL = `n4;    12'd281: toneL = `n4;    12'd282: toneL = `n4;    12'd283: toneL = `n4;    12'd284: toneL = `n4;    12'd285: toneL = `n4;    12'd286: toneL = `n4;    12'd287: toneL = `sil;    12'd288: toneL = `n5;    12'd289: toneL = `n5;    12'd290: toneL = `n5;    12'd291: toneL = `n5;    12'd292: toneL = `n5;    12'd293: toneL = `n5;    12'd294: toneL = `n5;    12'd295: toneL = `n5;    12'd296: toneL = `n5;    12'd297: toneL = `n5;    12'd298: toneL = `n5;    12'd299: toneL = `n5;    12'd300: toneL = `n5;    12'd301: toneL = `n5;    12'd302: toneL = `n5;    12'd303: toneL = `n5;    12'd304: toneL = `n5;    12'd305: toneL = `n5;    12'd306: toneL = `n5;    12'd307: toneL = `n5;    12'd308: toneL = `n5;    12'd309: toneL = `n5;    12'd310: toneL = `n5;    12'd311: toneL = `n5;    12'd312: toneL = `n5;    12'd313: toneL = `n5;    12'd314: toneL = `n5;    12'd315: toneL = `n5;    12'd316: toneL = `n5;    12'd317: toneL = `n5;    12'd318: toneL = `n5;    12'd319: toneL = `sil;
                12'd320: toneL = `n3;    12'd321: toneL = `n3;    12'd322: toneL = `n3;    12'd323: toneL = `n3;    12'd324: toneL = `n3;    12'd325: toneL = `n3;    12'd326: toneL = `n3;    12'd327: toneL = `n3;    12'd328: toneL = `n3;    12'd329: toneL = `n3;    12'd330: toneL = `n3;    12'd331: toneL = `n3;    12'd332: toneL = `n3;    12'd333: toneL = `n3;    12'd334: toneL = `n3;    12'd335: toneL = `sil;    12'd336: toneL = `n4;    12'd337: toneL = `n4;    12'd338: toneL = `n4;    12'd339: toneL = `n4;    12'd340: toneL = `n4;    12'd341: toneL = `n4;    12'd342: toneL = `n4;    12'd343: toneL = `n4;    12'd344: toneL = `n4;    12'd345: toneL = `n4;    12'd346: toneL = `n4;    12'd347: toneL = `n4;    12'd348: toneL = `n4;    12'd349: toneL = `n4;    12'd350: toneL = `n4;    12'd351: toneL = `sil;    12'd352: toneL = `n5;    12'd353: toneL = `n5;    12'd354: toneL = `n5;    12'd355: toneL = `n5;    12'd356: toneL = `n5;    12'd357: toneL = `n5;    12'd358: toneL = `n5;    12'd359: toneL = `n5;    12'd360: toneL = `n5;    12'd361: toneL = `n5;    12'd362: toneL = `n5;    12'd363: toneL = `n5;    12'd364: toneL = `n5;    12'd365: toneL = `n5;    12'd366: toneL = `n5;    12'd367: toneL = `n5;    12'd368: toneL = `n5;    12'd369: toneL = `n5;    12'd370: toneL = `n5;    12'd371: toneL = `n5;    12'd372: toneL = `n5;    12'd373: toneL = `n5;    12'd374: toneL = `n5;    12'd375: toneL = `n5;    12'd376: toneL = `n5;    12'd377: toneL = `n5;    12'd378: toneL = `n5;    12'd379: toneL = `n5;    12'd380: toneL = `n5;    12'd381: toneL = `n5;    12'd382: toneL = `n5;    12'd383: toneL = `sil;
                12'd384: toneL = `n5;    12'd385: toneL = `n5;    12'd386: toneL = `n5;    12'd387: toneL = `n5;    12'd388: toneL = `n5;    12'd389: toneL = `n5;    12'd390: toneL = `n5;    12'd391: toneL = `n5;    12'd392: toneL = `n5;    12'd393: toneL = `n5;    12'd394: toneL = `n5;    12'd395: toneL = `n5;    12'd396: toneL = `n5;    12'd397: toneL = `n5;    12'd398: toneL = `n5;    12'd399: toneL = `n5;    12'd400: toneL = `n5;    12'd401: toneL = `n5;    12'd402: toneL = `n5;    12'd403: toneL = `n5;    12'd404: toneL = `n5;    12'd405: toneL = `n5;    12'd406: toneL = `n5;    12'd407: toneL = `n5;    12'd408: toneL = `n5;    12'd409: toneL = `n5;    12'd410: toneL = `n5;    12'd411: toneL = `n5;    12'd412: toneL = `n5;    12'd413: toneL = `n5;    12'd414: toneL = `n5;    12'd415: toneL = `sil;    12'd416: toneL = `n3;    12'd417: toneL = `n3;    12'd418: toneL = `n3;    12'd419: toneL = `n3;    12'd420: toneL = `n3;    12'd421: toneL = `n3;    12'd422: toneL = `n3;    12'd423: toneL = `n3;    12'd424: toneL = `n3;    12'd425: toneL = `n3;    12'd426: toneL = `n3;    12'd427: toneL = `n3;    12'd428: toneL = `n3;    12'd429: toneL = `n3;    12'd430: toneL = `n3;    12'd431: toneL = `n3;    12'd432: toneL = `n3;    12'd433: toneL = `n3;    12'd434: toneL = `n3;    12'd435: toneL = `n3;    12'd436: toneL = `n3;    12'd437: toneL = `n3;    12'd438: toneL = `n3;    12'd439: toneL = `n3;    12'd440: toneL = `n3;    12'd441: toneL = `n3;    12'd442: toneL = `n3;    12'd443: toneL = `n3;    12'd444: toneL = `n3;    12'd445: toneL = `n3;    12'd446: toneL = `n3;    12'd447: toneL = `sil;
                12'd448: toneL = `n5;    12'd449: toneL = `n5;    12'd450: toneL = `n5;    12'd451: toneL = `n5;    12'd452: toneL = `n5;    12'd453: toneL = `n5;    12'd454: toneL = `n5;    12'd455: toneL = `n5;    12'd456: toneL = `n5;    12'd457: toneL = `n5;    12'd458: toneL = `n5;    12'd459: toneL = `n5;    12'd460: toneL = `n5;    12'd461: toneL = `n5;    12'd462: toneL = `n5;    12'd463: toneL = `n5;    12'd464: toneL = `n5;    12'd465: toneL = `n5;    12'd466: toneL = `n5;    12'd467: toneL = `n5;    12'd468: toneL = `n5;    12'd469: toneL = `n5;    12'd470: toneL = `n5;    12'd471: toneL = `n5;    12'd472: toneL = `n5;    12'd473: toneL = `n5;    12'd474: toneL = `n5;    12'd475: toneL = `n5;    12'd476: toneL = `n5;    12'd477: toneL = `n5;    12'd478: toneL = `n5;    12'd479: toneL = `sil;    12'd480: toneL = `n3;    12'd481: toneL = `n3;    12'd482: toneL = `n3;    12'd483: toneL = `n3;    12'd484: toneL = `n3;    12'd485: toneL = `n3;    12'd486: toneL = `n3;    12'd487: toneL = `n3;    12'd488: toneL = `n3;    12'd489: toneL = `n3;    12'd490: toneL = `n3;    12'd491: toneL = `n3;    12'd492: toneL = `n3;    12'd493: toneL = `n3;    12'd494: toneL = `n3;    12'd495: toneL = `n3;    12'd496: toneL = `n3;    12'd497: toneL = `n3;    12'd498: toneL = `n3;    12'd499: toneL = `n3;    12'd500: toneL = `n3;    12'd501: toneL = `n3;    12'd502: toneL = `n3;    12'd503: toneL = `n3;    12'd504: toneL = `n3;    12'd505: toneL = `n3;    12'd506: toneL = `n3;    12'd507: toneL = `n3;    12'd508: toneL = `n3;    12'd509: toneL = `n3;    12'd510: toneL = `n3;    12'd511: toneL = `sil;
                default : toneL = `sil;
            endcase
        end
        else begin
            toneL = `sil;
        end
    end
endmodule

//Jingle Bell
module music1 (
    input [11:0] ibeatNum,
    input en,
    output reg [31:0] toneL,
    output reg [31:0] toneR
);

    always @* begin
        if(en == 0) begin
            case(ibeatNum)
                12'd0: toneR = `s4;    12'd1: toneR = `s4;    12'd2: toneR = `s4;    12'd3: toneR = `s4;    12'd4: toneR = `s4;    12'd5: toneR = `s4;    12'd6: toneR = `s4;    12'd7: toneR = `sil;    12'd8: toneR = `s4;    12'd9: toneR = `s4;    12'd10: toneR = `s4;    12'd11: toneR = `s4;    12'd12: toneR = `s4;    12'd13: toneR = `s4;    12'd14: toneR = `s4;    12'd15: toneR = `sil;    12'd16: toneR = `s4;    12'd17: toneR = `s4;    12'd18: toneR = `s4;    12'd19: toneR = `s4;    12'd20: toneR = `s4;    12'd21: toneR = `s4;    12'd22: toneR = `s4;    12'd23: toneR = `s4;    12'd24: toneR = `s4;    12'd25: toneR = `s4;    12'd26: toneR = `s4;    12'd27: toneR = `s4;    12'd28: toneR = `s4;    12'd29: toneR = `s4;    12'd30: toneR = `s4;    12'd31: toneR = `sil;    12'd32: toneR = `s4;    12'd33: toneR = `s4;    12'd34: toneR = `s4;    12'd35: toneR = `s4;    12'd36: toneR = `s4;    12'd37: toneR = `s4;    12'd38: toneR = `s4;    12'd39: toneR = `sil;    12'd40: toneR = `s4;    12'd41: toneR = `s4;    12'd42: toneR = `s4;    12'd43: toneR = `s4;    12'd44: toneR = `s4;    12'd45: toneR = `s4;    12'd46: toneR = `s4;    12'd47: toneR = `sil;    12'd48: toneR = `s4;    12'd49: toneR = `s4;    12'd50: toneR = `s4;    12'd51: toneR = `s4;    12'd52: toneR = `s4;    12'd53: toneR = `s4;    12'd54: toneR = `s4;    12'd55: toneR = `s4;    12'd56: toneR = `s4;    12'd57: toneR = `s4;    12'd58: toneR = `s4;    12'd59: toneR = `s4;    12'd60: toneR = `s4;    12'd61: toneR = `s4;    12'd62: toneR = `s4;    12'd63: toneR = `sil;
                12'd64: toneR = `s4;    12'd65: toneR = `s4;    12'd66: toneR = `s4;    12'd67: toneR = `s4;    12'd68: toneR = `s4;    12'd69: toneR = `s4;    12'd70: toneR = `s4;    12'd71: toneR = `sil;    12'd72: toneR = `s6;    12'd73: toneR = `s6;    12'd74: toneR = `s6;    12'd75: toneR = `s6;    12'd76: toneR = `s6;    12'd77: toneR = `s6;    12'd78: toneR = `s6;    12'd79: toneR = `sil;    12'd80: toneR = `s2;    12'd81: toneR = `s2;    12'd82: toneR = `s2;    12'd83: toneR = `s2;    12'd84: toneR = `s2;    12'd85: toneR = `s2;    12'd86: toneR = `s2;    12'd87: toneR = `s2;    12'd88: toneR = `s2;    12'd89: toneR = `s2;    12'd90: toneR = `s2;    12'd91: toneR = `sil;    12'd92: toneR = `s3;    12'd93: toneR = `s3;    12'd94: toneR = `s3;    12'd95: toneR = `sil;    12'd96: toneR = `s4;    12'd97: toneR = `s4;    12'd98: toneR = `s4;    12'd99: toneR = `s4;    12'd100: toneR = `s4;    12'd101: toneR = `s4;    12'd102: toneR = `s4;    12'd103: toneR = `s4;    12'd104: toneR = `s4;    12'd105: toneR = `s4;    12'd106: toneR = `s4;    12'd107: toneR = `s4;    12'd108: toneR = `s4;    12'd109: toneR = `s4;    12'd110: toneR = `s4;    12'd111: toneR = `s4;    12'd112: toneR = `s4;    12'd113: toneR = `s4;    12'd114: toneR = `s4;    12'd115: toneR = `s4;    12'd116: toneR = `s4;    12'd117: toneR = `s4;    12'd118: toneR = `s4;    12'd119: toneR = `s4;    12'd120: toneR = `s4;    12'd121: toneR = `s4;    12'd122: toneR = `s4;    12'd123: toneR = `s4;    12'd124: toneR = `s4;    12'd125: toneR = `s4;    12'd126: toneR = `s4;    12'd127: toneR = `sil;
                12'd128: toneR = `s5;    12'd129: toneR = `s5;    12'd130: toneR = `s5;    12'd131: toneR = `s5;    12'd132: toneR = `s5;    12'd133: toneR = `s5;    12'd134: toneR = `s5;    12'd135: toneR = `sil;    12'd136: toneR = `s5;    12'd137: toneR = `s5;    12'd138: toneR = `s5;    12'd139: toneR = `s5;    12'd140: toneR = `s5;    12'd141: toneR = `s5;    12'd142: toneR = `s5;    12'd143: toneR = `sil;    12'd144: toneR = `s5;    12'd145: toneR = `s5;    12'd146: toneR = `s5;    12'd147: toneR = `s5;    12'd148: toneR = `s5;    12'd149: toneR = `s5;    12'd150: toneR = `s5;    12'd151: toneR = `s5;    12'd152: toneR = `s5;    12'd153: toneR = `s5;    12'd154: toneR = `s5;    12'd155: toneR = `sil;    12'd156: toneR = `s5;    12'd157: toneR = `s5;    12'd158: toneR = `s5;    12'd187: toneR = `sil;    12'd160: toneR = `s5;    12'd161: toneR = `s5;    12'd162: toneR = `s5;    12'd163: toneR = `s5;    12'd164: toneR = `s5;    12'd165: toneR = `s5;    12'd166: toneR = `s5;    12'd167: toneR = `sil;    12'd168: toneR = `s4;    12'd169: toneR = `s4;    12'd170: toneR = `s4;    12'd171: toneR = `s4;    12'd172: toneR = `s4;    12'd173: toneR = `s4;    12'd174: toneR = `s4;    12'd175: toneR = `sil;    12'd176: toneR = `s4;    12'd177: toneR = `s4;    12'd178: toneR = `s4;    12'd179: toneR = `s4;    12'd180: toneR = `s4;    12'd181: toneR = `s4;    12'd182: toneR = `s4;    12'd183: toneR = `s4;    12'd184: toneR = `s4;    12'd185: toneR = `s4;    12'd186: toneR = `s4;    12'd187: toneR = `s4;    12'd188: toneR = `s4;    12'd189: toneR = `s4;    12'd190: toneR = `s4;    12'd191: toneR = `sil;
                12'd192: toneR = `s4;    12'd193: toneR = `s4;    12'd194: toneR = `s4;    12'd195: toneR = `s4;    12'd196: toneR = `s4;    12'd197: toneR = `s4;    12'd198: toneR = `s4;    12'd199: toneR = `sil;    12'd200: toneR = `s3;    12'd201: toneR = `s3;    12'd202: toneR = `s3;    12'd203: toneR = `s3;    12'd204: toneR = `s3;    12'd205: toneR = `s3;    12'd206: toneR = `s3;    12'd207: toneR = `sil;    12'd208: toneR = `s3;    12'd209: toneR = `s3;    12'd210: toneR = `s3;    12'd211: toneR = `s3;    12'd212: toneR = `s3;    12'd213: toneR = `s3;    12'd214: toneR = `s3;    12'd215: toneR = `sil;    12'd216: toneR = `s4;    12'd217: toneR = `s4;    12'd218: toneR = `s4;    12'd219: toneR = `s4;    12'd220: toneR = `s4;    12'd221: toneR = `s4;    12'd222: toneR = `s4;    12'd223: toneR = `sil;    12'd224: toneR = `s3;    12'd225: toneR = `s3;    12'd226: toneR = `s3;    12'd227: toneR = `s3;    12'd228: toneR = `s3;    12'd229: toneR = `s3;    12'd230: toneR = `s3;    12'd231: toneR = `s3;    12'd232: toneR = `s3;    12'd233: toneR = `s3;    12'd234: toneR = `s3;    12'd235: toneR = `s3;    12'd236: toneR = `s3;    12'd237: toneR = `s3;    12'd238: toneR = `s3;    12'd239: toneR = `sil;    12'd240: toneR = `s6;    12'd241: toneR = `s6;    12'd242: toneR = `s6;    12'd243: toneR = `s6;    12'd244: toneR = `s6;    12'd245: toneR = `s6;    12'd246: toneR = `s6;    12'd247: toneR = `s6;    12'd248: toneR = `s6;    12'd249: toneR = `s6;    12'd250: toneR = `s6;    12'd251: toneR = `s6;    12'd252: toneR = `s6;    12'd253: toneR = `s6;    12'd254: toneR = `s6;    12'd255: toneR = `sil;
                12'd256: toneR = `s4;    12'd257: toneR = `s4;    12'd258: toneR = `s4;    12'd259: toneR = `s4;    12'd260: toneR = `s4;    12'd261: toneR = `s4;    12'd262: toneR = `s4;    12'd263: toneR = `sil;    12'd264: toneR = `s4;    12'd265: toneR = `s4;    12'd266: toneR = `s4;    12'd267: toneR = `s4;    12'd268: toneR = `s4;    12'd269: toneR = `s4;    12'd270: toneR = `s4;    12'd271: toneR = `sil;    12'd272: toneR = `s4;    12'd273: toneR = `s4;    12'd274: toneR = `s4;    12'd275: toneR = `s4;    12'd276: toneR = `s4;    12'd277: toneR = `s4;    12'd278: toneR = `s4;    12'd279: toneR = `s4;    12'd280: toneR = `s4;    12'd281: toneR = `s4;    12'd282: toneR = `s4;    12'd283: toneR = `s4;    12'd284: toneR = `s4;    12'd285: toneR = `s4;    12'd286: toneR = `s4;    12'd287: toneR = `sil;    12'd288: toneR = `s4;    12'd289: toneR = `s4;    12'd290: toneR = `s4;    12'd291: toneR = `s4;    12'd292: toneR = `s4;    12'd293: toneR = `s4;    12'd294: toneR = `s4;    12'd295: toneR = `sil;    12'd296: toneR = `s4;    12'd297: toneR = `s4;    12'd298: toneR = `s4;    12'd299: toneR = `s4;    12'd300: toneR = `s4;    12'd301: toneR = `s4;    12'd302: toneR = `s4;    12'd303: toneR = `sil;    12'd304: toneR = `s4;    12'd305: toneR = `s4;    12'd306: toneR = `s4;    12'd307: toneR = `s4;    12'd308: toneR = `s4;    12'd309: toneR = `s4;    12'd310: toneR = `s4;    12'd311: toneR = `s4;    12'd312: toneR = `s4;    12'd313: toneR = `s4;    12'd314: toneR = `s4;    12'd315: toneR = `s4;    12'd316: toneR = `s4;    12'd317: toneR = `s4;    12'd318: toneR = `s4;    12'd319: toneR = `sil;
                12'd320: toneR = `s4;    12'd321: toneR = `s4;    12'd322: toneR = `s4;    12'd323: toneR = `s4;    12'd324: toneR = `s4;    12'd325: toneR = `s4;    12'd326: toneR = `s4;    12'd327: toneR = `sil;    12'd328: toneR = `s6;    12'd329: toneR = `s6;    12'd330: toneR = `s6;    12'd331: toneR = `s6;    12'd332: toneR = `s6;    12'd333: toneR = `s6;    12'd334: toneR = `s6;    12'd335: toneR = `sil;    12'd336: toneR = `s2;    12'd337: toneR = `s2;    12'd338: toneR = `s2;    12'd339: toneR = `s2;    12'd340: toneR = `s2;    12'd341: toneR = `s2;    12'd342: toneR = `s2;    12'd343: toneR = `s2;    12'd344: toneR = `s2;    12'd345: toneR = `s2;    12'd346: toneR = `s2;    12'd347: toneR = `sil;    12'd348: toneR = `s3;    12'd349: toneR = `s3;    12'd350: toneR = `s3;    12'd351: toneR = `sil;    12'd352: toneR = `s4;    12'd353: toneR = `s4;    12'd354: toneR = `s4;    12'd355: toneR = `s4;    12'd356: toneR = `s4;    12'd357: toneR = `s4;    12'd358: toneR = `s4;    12'd359: toneR = `s4;    12'd360: toneR = `s4;    12'd361: toneR = `s4;    12'd362: toneR = `s4;    12'd363: toneR = `s4;    12'd364: toneR = `s4;    12'd365: toneR = `s4;    12'd366: toneR = `s4;    12'd367: toneR = `s4;    12'd368: toneR = `s4;    12'd369: toneR = `s4;    12'd370: toneR = `s4;    12'd371: toneR = `s4;    12'd372: toneR = `s4;    12'd373: toneR = `s4;    12'd374: toneR = `s4;    12'd375: toneR = `s4;    12'd376: toneR = `s4;    12'd377: toneR = `s4;    12'd378: toneR = `s4;    12'd379: toneR = `s4;    12'd380: toneR = `s4;    12'd381: toneR = `s4;    12'd382: toneR = `s4;    12'd383: toneR = `sil;
                12'd384: toneR = `s5;    12'd385: toneR = `s5;    12'd386: toneR = `s5;    12'd387: toneR = `s5;    12'd388: toneR = `s5;    12'd389: toneR = `s5;    12'd390: toneR = `s5;    12'd391: toneR = `sil;    12'd392: toneR = `s5;    12'd393: toneR = `s5;    12'd394: toneR = `s5;    12'd395: toneR = `s5;    12'd396: toneR = `s5;    12'd397: toneR = `s5;    12'd398: toneR = `s5;    12'd399: toneR = `sil;    12'd400: toneR = `s5;    12'd401: toneR = `s5;    12'd402: toneR = `s5;    12'd403: toneR = `s5;    12'd404: toneR = `s5;    12'd405: toneR = `s5;    12'd406: toneR = `s5;    12'd407: toneR = `s5;    12'd408: toneR = `s5;    12'd409: toneR = `s5;    12'd410: toneR = `s5;    12'd411: toneR = `sil;    12'd412: toneR = `s5;    12'd413: toneR = `s5;    12'd414: toneR = `s5;    12'd415: toneR = `sil;    12'd416: toneR = `s5;    12'd417: toneR = `s5;    12'd418: toneR = `s5;    12'd419: toneR = `s5;    12'd420: toneR = `s5;    12'd421: toneR = `s5;    12'd422: toneR = `s5;    12'd423: toneR = `sil;    12'd424: toneR = `s4;    12'd425: toneR = `s4;    12'd426: toneR = `s4;    12'd427: toneR = `s4;    12'd428: toneR = `s4;    12'd429: toneR = `s4;    12'd430: toneR = `s4;    12'd431: toneR = `sil;    12'd432: toneR = `s5;    12'd433: toneR = `s5;    12'd434: toneR = `s5;    12'd435: toneR = `s5;    12'd436: toneR = `s5;    12'd437: toneR = `s5;    12'd438: toneR = `s5;    12'd439: toneR = `s5;    12'd440: toneR = `s5;    12'd441: toneR = `s5;    12'd442: toneR = `s5;    12'd443: toneR = `s5;    12'd444: toneR = `s5;    12'd445: toneR = `s5;    12'd446: toneR = `s5;    12'd447: toneR = `sil;
                12'd448: toneR = `s6;    12'd449: toneR = `s6;    12'd450: toneR = `s6;    12'd451: toneR = `s6;    12'd452: toneR = `s6;    12'd453: toneR = `s6;    12'd454: toneR = `s6;    12'd455: toneR = `sil;    12'd456: toneR = `s6;    12'd457: toneR = `s6;    12'd458: toneR = `s6;    12'd459: toneR = `s6;    12'd460: toneR = `s6;    12'd461: toneR = `s6;    12'd462: toneR = `s6;    12'd463: toneR = `sil;    12'd464: toneR = `s5;    12'd465: toneR = `s5;    12'd466: toneR = `s5;    12'd467: toneR = `s5;    12'd468: toneR = `s5;    12'd469: toneR = `s5;    12'd470: toneR = `s5;    12'd471: toneR = `sil;    12'd472: toneR = `s3;    12'd473: toneR = `s3;    12'd474: toneR = `s3;    12'd475: toneR = `s3;    12'd476: toneR = `s3;    12'd477: toneR = `s3;    12'd478: toneR = `s3;    12'd479: toneR = `sil;    12'd480: toneR = `s2;    12'd481: toneR = `s2;    12'd482: toneR = `s2;    12'd483: toneR = `s2;    12'd484: toneR = `s2;    12'd485: toneR = `s2;    12'd486: toneR = `s2;    12'd487: toneR = `s2;    12'd488: toneR = `s2;    12'd489: toneR = `s2;    12'd490: toneR = `s2;    12'd491: toneR = `s2;    12'd492: toneR = `s2;    12'd493: toneR = `s2;    12'd494: toneR = `s2;    12'd495: toneR = `s2;    12'd496: toneR = `s2;    12'd497: toneR = `s2;    12'd498: toneR = `s2;    12'd499: toneR = `s2;    12'd500: toneR = `s2;    12'd501: toneR = `s2;    12'd502: toneR = `s2;    12'd503: toneR = `s2;    12'd504: toneR = `s2;    12'd505: toneR = `s2;    12'd506: toneR = `s2;    12'd507: toneR = `s2;    12'd508: toneR = `s2;    12'd509: toneR = `s2;    12'd510: toneR = `s2;    12'd511: toneR = `sil;
                default : toneR = `sil;
            endcase
        end else begin
            toneR = `sil;
        end
    end

    always @(*) begin
        if(en==0)begin
            case(ibeatNum)
                12'd0: toneL = `n2;    12'd1: toneL = `n2;    12'd2: toneL = `n2;    12'd3: toneL = `n2;    12'd4: toneL = `n2;    12'd5: toneL = `n2;    12'd6: toneL = `n2;    12'd7: toneL = `n2;    12'd8: toneL = `n6;    12'd9: toneL = `n6;    12'd10: toneL = `n6;    12'd11: toneL = `n6;    12'd12: toneL = `n6;    12'd13: toneL = `n6;    12'd14: toneL = `n6;    12'd15: toneL = `n6;    12'd16: toneL = `n4;    12'd17: toneL = `n4;    12'd18: toneL = `n4;    12'd19: toneL = `n4;    12'd20: toneL = `n4;    12'd21: toneL = `n4;    12'd22: toneL = `n4;    12'd23: toneL = `n4;    12'd24: toneL = `n6;    12'd25: toneL = `n6;    12'd26: toneL = `n6;    12'd27: toneL = `n6;    12'd28: toneL = `n6;    12'd29: toneL = `n6;    12'd30: toneL = `n6;    12'd31: toneL = `sil;    12'd32: toneL = `n2;    12'd33: toneL = `n2;    12'd34: toneL = `n2;    12'd35: toneL = `n2;    12'd36: toneL = `n2;    12'd37: toneL = `n2;    12'd38: toneL = `n2;    12'd39: toneL = `n2;    12'd40: toneL = `n6;    12'd41: toneL = `n6;    12'd42: toneL = `n6;    12'd43: toneL = `n6;    12'd44: toneL = `n6;    12'd45: toneL = `n6;    12'd46: toneL = `n6;    12'd47: toneL = `n6;    12'd48: toneL = `n4;    12'd49: toneL = `n4;    12'd50: toneL = `n4;    12'd51: toneL = `n4;    12'd52: toneL = `n4;    12'd53: toneL = `n4;    12'd54: toneL = `n4;    12'd55: toneL = `n4;    12'd56: toneL = `n6;    12'd57: toneL = `n6;    12'd58: toneL = `n6;    12'd59: toneL = `n6;    12'd60: toneL = `n6;    12'd61: toneL = `n6;    12'd62: toneL = `n6;    12'd63: toneL = `sil;
                12'd64: toneL = `n2;    12'd65: toneL = `n2;    12'd66: toneL = `n2;    12'd67: toneL = `n2;    12'd68: toneL = `n2;    12'd69: toneL = `n2;    12'd70: toneL = `n2;    12'd71: toneL = `n2;    12'd72: toneL = `n6;    12'd73: toneL = `n6;    12'd74: toneL = `n6;    12'd75: toneL = `n6;    12'd76: toneL = `n6;    12'd77: toneL = `n6;    12'd78: toneL = `n6;    12'd79: toneL = `n6;    12'd80: toneL = `n4;    12'd81: toneL = `n4;    12'd82: toneL = `n4;    12'd83: toneL = `n4;    12'd84: toneL = `n4;    12'd85: toneL = `n4;    12'd86: toneL = `n4;    12'd87: toneL = `n4;    12'd88: toneL = `n6;    12'd89: toneL = `n6;    12'd90: toneL = `n6;    12'd91: toneL = `n6;    12'd92: toneL = `n6;    12'd93: toneL = `n6;    12'd94: toneL = `n6;    12'd95: toneL = `sil;    12'd96: toneL = `n2;    12'd97: toneL = `n2;    12'd98: toneL = `n2;    12'd99: toneL = `n2;    12'd100: toneL = `n2;    12'd101: toneL = `n2;    12'd102: toneL = `n2;    12'd103: toneL = `n2;    12'd104: toneL = `n6;    12'd105: toneL = `n6;    12'd106: toneL = `n6;    12'd107: toneL = `n6;    12'd108: toneL = `n6;    12'd109: toneL = `n6;    12'd110: toneL = `n6;    12'd111: toneL = `n6;    12'd112: toneL = `n4;    12'd113: toneL = `n4;    12'd114: toneL = `n4;    12'd115: toneL = `n4;    12'd116: toneL = `n4;    12'd117: toneL = `n4;    12'd118: toneL = `n4;    12'd119: toneL = `n4;    12'd120: toneL = `n6;    12'd121: toneL = `n6;    12'd122: toneL = `n6;    12'd123: toneL = `n6;    12'd124: toneL = `n6;    12'd125: toneL = `n6;    12'd126: toneL = `n6;    12'd127: toneL = `sil;
                12'd128: toneL = `n2;    12'd129: toneL = `n2;    12'd130: toneL = `n2;    12'd131: toneL = `n2;    12'd132: toneL = `n2;    12'd133: toneL = `n2;    12'd134: toneL = `n2;    12'd135: toneL = `n2;    12'd136: toneL = `n7;    12'd137: toneL = `n7;    12'd138: toneL = `n7;    12'd139: toneL = `n7;    12'd140: toneL = `n7;    12'd141: toneL = `n7;    12'd142: toneL = `n7;    12'd143: toneL = `n7;    12'd144: toneL = `n5;    12'd145: toneL = `n5;    12'd146: toneL = `n5;    12'd147: toneL = `n5;    12'd148: toneL = `n5;    12'd149: toneL = `n5;    12'd150: toneL = `n5;    12'd151: toneL = `n5;    12'd152: toneL = `n7;    12'd153: toneL = `n7;    12'd154: toneL = `n7;    12'd155: toneL = `n7;    12'd156: toneL = `n7;    12'd157: toneL = `n7;    12'd158: toneL = `n7;    12'd159: toneL = `sil;    12'd160: toneL = `n2;    12'd161: toneL = `n2;    12'd162: toneL = `n2;    12'd163: toneL = `n2;    12'd164: toneL = `n2;    12'd165: toneL = `n2;    12'd166: toneL = `n2;    12'd167: toneL = `n2;    12'd168: toneL = `n6;    12'd169: toneL = `n6;    12'd170: toneL = `n6;    12'd171: toneL = `n6;    12'd172: toneL = `n6;    12'd173: toneL = `n6;    12'd174: toneL = `n6;    12'd175: toneL = `n6;    12'd176: toneL = `n4;    12'd177: toneL = `n4;    12'd178: toneL = `n4;    12'd179: toneL = `n4;    12'd180: toneL = `n4;    12'd181: toneL = `n4;    12'd182: toneL = `n4;    12'd183: toneL = `n4;    12'd184: toneL = `n6;    12'd185: toneL = `n6;    12'd186: toneL = `n6;    12'd187: toneL = `n6;    12'd188: toneL = `n6;    12'd189: toneL = `n6;    12'd190: toneL = `n6;    12'd191: toneL = `sil;
                12'd192: toneL = `n6;    12'd193: toneL = `n6;    12'd194: toneL = `n6;    12'd195: toneL = `n6;    12'd196: toneL = `n6;    12'd197: toneL = `n6;    12'd198: toneL = `n6;    12'd199: toneL = `n6;    12'd200: toneL = `n6;    12'd201: toneL = `n6;    12'd202: toneL = `n6;    12'd203: toneL = `n6;    12'd204: toneL = `n6;    12'd205: toneL = `n6;    12'd206: toneL = `n6;    12'd207: toneL = `sil;    12'd208: toneL = `n3;    12'd209: toneL = `n3;    12'd210: toneL = `n3;    12'd211: toneL = `n3;    12'd212: toneL = `n3;    12'd213: toneL = `n3;    12'd214: toneL = `n3;    12'd215: toneL = `n3;    12'd216: toneL = `n3;    12'd217: toneL = `n3;    12'd218: toneL = `n3;    12'd219: toneL = `n3;    12'd220: toneL = `n3;    12'd221: toneL = `n3;    12'd222: toneL = `n3;    12'd223: toneL = `sil;    12'd224: toneL = `n6;    12'd225: toneL = `n6;    12'd226: toneL = `n6;    12'd227: toneL = `n6;    12'd228: toneL = `n6;    12'd229: toneL = `n6;    12'd230: toneL = `n6;    12'd231: toneL = `n6;    12'd232: toneL = `n5;    12'd233: toneL = `n5;    12'd234: toneL = `n5;    12'd235: toneL = `n5;    12'd236: toneL = `n5;    12'd237: toneL = `n5;    12'd238: toneL = `n5;    12'd239: toneL = `n5;    12'd240: toneL = `n4;    12'd241: toneL = `n4;    12'd242: toneL = `n4;    12'd243: toneL = `n4;    12'd244: toneL = `n4;    12'd245: toneL = `n4;    12'd246: toneL = `n4;    12'd247: toneL = `sil;    12'd248: toneL = `n4;    12'd249: toneL = `n4;    12'd250: toneL = `n4;    12'd251: toneL = `n4;    12'd252: toneL = `n4;    12'd253: toneL = `n4;    12'd254: toneL = `n4;    12'd255: toneL = `sil;
                12'd256: toneL = `n4;    12'd257: toneL = `n4;    12'd258: toneL = `n4;    12'd259: toneL = `n4;    12'd260: toneL = `n4;    12'd261: toneL = `n4;    12'd262: toneL = `n4;    12'd263: toneL = `n4;    12'd264: toneL = `n6;    12'd265: toneL = `n6;    12'd266: toneL = `n6;    12'd267: toneL = `n6;    12'd268: toneL = `n6;    12'd269: toneL = `n6;    12'd270: toneL = `n6;    12'd271: toneL = `n6;    12'd272: toneL = `n4;    12'd273: toneL = `n4;    12'd274: toneL = `n4;    12'd275: toneL = `n4;    12'd276: toneL = `n4;    12'd277: toneL = `n4;    12'd278: toneL = `n4;    12'd279: toneL = `n4;    12'd280: toneL = `n6;    12'd281: toneL = `n6;    12'd282: toneL = `n6;    12'd283: toneL = `n6;    12'd284: toneL = `n6;    12'd285: toneL = `n6;    12'd286: toneL = `n6;    12'd287: toneL = `sil;    12'd288: toneL = `n2;    12'd289: toneL = `n2;    12'd290: toneL = `n2;    12'd291: toneL = `n2;    12'd292: toneL = `n2;    12'd293: toneL = `n2;    12'd294: toneL = `n2;    12'd295: toneL = `n2;    12'd296: toneL = `n6;    12'd297: toneL = `n6;    12'd298: toneL = `n6;    12'd299: toneL = `n6;    12'd300: toneL = `n6;    12'd301: toneL = `n6;    12'd302: toneL = `n6;    12'd303: toneL = `n6;    12'd304: toneL = `n4;    12'd305: toneL = `n4;    12'd306: toneL = `n4;    12'd307: toneL = `n4;    12'd308: toneL = `n4;    12'd309: toneL = `n4;    12'd310: toneL = `n4;    12'd311: toneL = `n4;    12'd312: toneL = `n6;    12'd313: toneL = `n6;    12'd314: toneL = `n6;    12'd315: toneL = `n6;    12'd316: toneL = `n6;    12'd317: toneL = `n6;    12'd318: toneL = `n6;    12'd319: toneL = `sil;
                12'd320: toneL = `n2;    12'd321: toneL = `n2;    12'd322: toneL = `n2;    12'd323: toneL = `n2;    12'd324: toneL = `n2;    12'd325: toneL = `n2;    12'd326: toneL = `n2;    12'd327: toneL = `n2;    12'd328: toneL = `n6;    12'd329: toneL = `n6;    12'd330: toneL = `n6;    12'd331: toneL = `n6;    12'd332: toneL = `n6;    12'd333: toneL = `n6;    12'd334: toneL = `n6;    12'd335: toneL = `n6;    12'd336: toneL = `n4;    12'd337: toneL = `n4;    12'd338: toneL = `n4;    12'd339: toneL = `n4;    12'd340: toneL = `n4;    12'd341: toneL = `n4;    12'd342: toneL = `n4;    12'd343: toneL = `n4;    12'd344: toneL = `n6;    12'd345: toneL = `n6;    12'd346: toneL = `n6;    12'd347: toneL = `n6;    12'd348: toneL = `n6;    12'd349: toneL = `n6;    12'd350: toneL = `n6;    12'd351: toneL = `sil;    12'd352: toneL = `n2;    12'd353: toneL = `n2;    12'd354: toneL = `n2;    12'd355: toneL = `n2;    12'd356: toneL = `n2;    12'd357: toneL = `n2;    12'd358: toneL = `n2;    12'd359: toneL = `n2;    12'd360: toneL = `n6;    12'd361: toneL = `n6;    12'd362: toneL = `n6;    12'd363: toneL = `n6;    12'd364: toneL = `n6;    12'd365: toneL = `n6;    12'd366: toneL = `n6;    12'd367: toneL = `n6;    12'd368: toneL = `n4;    12'd369: toneL = `n4;    12'd370: toneL = `n4;    12'd371: toneL = `n4;    12'd372: toneL = `n4;    12'd373: toneL = `n4;    12'd374: toneL = `n4;    12'd375: toneL = `n4;    12'd376: toneL = `n6;    12'd377: toneL = `n6;    12'd378: toneL = `n6;    12'd379: toneL = `n6;    12'd380: toneL = `n6;    12'd381: toneL = `n6;    12'd382: toneL = `n6;    12'd383: toneL = `sil;
                12'd384: toneL = `n2;    12'd385: toneL = `n2;    12'd386: toneL = `n2;    12'd387: toneL = `n2;    12'd388: toneL = `n2;    12'd389: toneL = `n2;    12'd390: toneL = `n2;    12'd391: toneL = `n2;    12'd392: toneL = `n7;    12'd393: toneL = `n7;    12'd394: toneL = `n7;    12'd395: toneL = `n7;    12'd396: toneL = `n7;    12'd397: toneL = `n7;    12'd398: toneL = `n7;    12'd399: toneL = `n7;    12'd400: toneL = `n5;    12'd401: toneL = `n5;    12'd402: toneL = `n5;    12'd403: toneL = `n5;    12'd404: toneL = `n5;    12'd405: toneL = `n5;    12'd406: toneL = `n5;    12'd407: toneL = `n5;    12'd408: toneL = `n7;    12'd409: toneL = `n7;    12'd410: toneL = `n7;    12'd411: toneL = `n7;    12'd412: toneL = `n7;    12'd413: toneL = `n7;    12'd414: toneL = `n7;    12'd415: toneL = `sil;    12'd416: toneL = `n2;    12'd417: toneL = `n2;    12'd418: toneL = `n2;    12'd419: toneL = `n2;    12'd420: toneL = `n2;    12'd421: toneL = `n2;    12'd422: toneL = `n2;    12'd423: toneL = `n2;    12'd424: toneL = `n6;    12'd425: toneL = `n6;    12'd426: toneL = `n6;    12'd427: toneL = `n6;    12'd428: toneL = `n6;    12'd429: toneL = `n6;    12'd430: toneL = `n6;    12'd431: toneL = `n6;    12'd432: toneL = `n4;    12'd433: toneL = `n4;    12'd434: toneL = `n4;    12'd435: toneL = `n4;    12'd436: toneL = `n4;    12'd437: toneL = `n4;    12'd438: toneL = `n4;    12'd439: toneL = `n4;    12'd440: toneL = `n6;    12'd441: toneL = `n6;    12'd442: toneL = `n6;    12'd443: toneL = `n6;    12'd444: toneL = `n6;    12'd445: toneL = `n6;    12'd446: toneL = `n6;    12'd447: toneL = `sil;
                12'd448: toneL = `n2;    12'd449: toneL = `n2;    12'd450: toneL = `n2;    12'd451: toneL = `n2;    12'd452: toneL = `n2;    12'd453: toneL = `n2;    12'd454: toneL = `n2;    12'd455: toneL = `n2;    12'd456: toneL = `n6;    12'd457: toneL = `n6;    12'd458: toneL = `n6;    12'd459: toneL = `n6;    12'd460: toneL = `n6;    12'd461: toneL = `n6;    12'd462: toneL = `n6;    12'd463: toneL = `n6;    12'd464: toneL = `s1;    12'd465: toneL = `s1;    12'd466: toneL = `s1;    12'd467: toneL = `s1;    12'd468: toneL = `s1;    12'd469: toneL = `s1;    12'd470: toneL = `s1;    12'd471: toneL = `s1;    12'd472: toneL = `n6;    12'd473: toneL = `n6;    12'd474: toneL = `n6;    12'd475: toneL = `n6;    12'd476: toneL = `n6;    12'd477: toneL = `n6;    12'd478: toneL = `n6;    12'd479: toneL = `sil;    12'd480: toneL = `s2;    12'd481: toneL = `s2;    12'd482: toneL = `s2;    12'd483: toneL = `s2;    12'd484: toneL = `s2;    12'd485: toneL = `s2;    12'd486: toneL = `s2;    12'd487: toneL = `s2;    12'd488: toneL = `n6;    12'd489: toneL = `n6;    12'd490: toneL = `n6;    12'd491: toneL = `n6;    12'd492: toneL = `n6;    12'd493: toneL = `n6;    12'd494: toneL = `n6;    12'd495: toneL = `sil;    12'd496: toneL = `n2;    12'd497: toneL = `n2;    12'd498: toneL = `n2;    12'd499: toneL = `n2;    12'd500: toneL = `n2;    12'd501: toneL = `n2;    12'd502: toneL = `n2;    12'd503: toneL = `n2;    12'd504: toneL = `n2;    12'd505: toneL = `n2;    12'd506: toneL = `n2;    12'd507: toneL = `n2;    12'd508: toneL = `n2;    12'd509: toneL = `n2;    12'd510: toneL = `n2;    12'd511: toneL = `sil;
                default : toneL = `sil;
            endcase
        end
        else begin
            toneL = `sil;
        end
    end
endmodule